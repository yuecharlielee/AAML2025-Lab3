module PE(
    
);
endmodule